library verilog;
use verilog.vl_types.all;
entity Digtal_Main_vlg_tst is
end Digtal_Main_vlg_tst;
